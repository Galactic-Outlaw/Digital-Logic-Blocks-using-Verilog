module clock(y,x);
input x;
output y;
not n1(y,x);
endmodule