module mux8_1_if_testmodule();
reg [7:0] D;
reg [2:0] S;
wire P;
mux8_1_if test(P,D,S);
initial
begin
$dumpfile("mux8_1_if_test.vcd");
$dumpvars(0,mux8_1_if_testmodule);
end
initial
begin
D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=0;
S[0]=0;
S[1]=0;
S[2]=0;
#10;

D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=1;
D[5]=0;
D[6]=1;
D[7]=1;
S[0]=0;
S[1]=0;
S[2]=1;
#10;

D[0]=0;
D[1]=0;
D[2]=0;
D[3]=1;
D[4]=1;
D[5]=1;
D[6]=0;
D[7]=0;
S[0]=0;
S[1]=1;
S[2]=0;
#10;

D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=1;
D[5]=0;
D[6]=1;
D[7]=0;
S[0]=0;
S[1]=1;
S[2]=1;
#10;

D[0]=0;
D[1]=0;
D[2]=0;
D[3]=1;
D[4]=0;
D[5]=1;
D[6]=0;
D[7]=0;
S[0]=1;
S[1]=0;
S[2]=0;
#10;

D[0]=0;
D[1]=0;
D[2]=0;
D[3]=1;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=1;
S[0]=1;
S[1]=0;
S[2]=1;
#10;

D[0]=0;
D[1]=0;
D[2]=0;
D[3]=1;
D[4]=0;
D[5]=0;
D[6]=1;
D[7]=0;
S[0]=1;
S[1]=1;
S[2]=0;
#10;

D[0]=1;
D[1]=1;
D[2]=1;
D[3]=1;
D[4]=1;
D[5]=1;
D[6]=1;
D[7]=1;
S[0]=1;
S[1]=1;
S[2]=1;
#10;


end
endmodule
