module mux8to3_en_testmodule();
reg [7:0] D;
wire [2:0] Q;
mux8to3_en test (Q,D);
initial
begin
$dumpfile("mux8to3_en_test.vcd");
$dumpvars(0,mux8to3_en_testmodule);
end
initial
begin
D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=0;
#10;
D[0]=1;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=0;
#10;
D[0]=0;
D[1]=1;
D[2]=0;
D[3]=0;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=0;
#10;
D[0]=0;
D[1]=0;
D[2]=1;
D[3]=0;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=0;
#10;
D[0]=0;
D[1]=0;
D[2]=0;
D[3]=1;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=0;
#10;
D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=1;
D[5]=0;
D[6]=0;
D[7]=0;
#10;
D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=0;
D[5]=1;
D[6]=0;
D[7]=0;
#10;
D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=0;
D[5]=0;
D[6]=1;
D[7]=0;
#10;
D[0]=0;
D[1]=0;
D[2]=0;
D[3]=0;
D[4]=0;
D[5]=0;
D[6]=0;
D[7]=1;
#10;
end
endmodule